//??????????
module AddBranch#(parameter WIDTH=32)(inAddr_add,inAddr_sl2,outAddr);
  input[WIDTH-1:0] inAddr_add;//??pc?4???????
  input[WIDTH-1:0] inAddr_sl2;//??????????
  output[WIDTH-1:0] outAddr;
  
  assign outAddr=inAddr_add+inAddr_sl2;
   
endmodule
